library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      endereco : in  unsigned(7 downto 0);
      dado     : out unsigned(18 downto 0)
   );
end entity;

architecture a_rom of rom is
   type mem is array (0 to 255) of unsigned(18 downto 0);

   constant conteudo_rom : mem := (
      ---- *****PASSO 1: colocar os valores de 1 a 32 ****** ----

      ---- SETUP INICIAL ----
      0  => "1001" & "000" & "000" & "100000001",  -- LD ACC,#1
      
      1  => "1111" & "001" & "000" & "000000001",  -- MOV R1,ACC

      2  => "1001" & "000" & "000" & "000100000",  -- ACC = 32
      
      3  => "1111" & "010" & "000" & "000000000",  -- R2 = 32
      
      -- INICIO DO LOOP
      4  => "1001" & "000" & "000" & "000000000",  -- ACC = 0

      5  => "1111" & "011" & "000" & "000000000",  -- MOV, R3, ACC

      6  => "0110" & "001" & "000" & "000000000",  -- ADD, R1, ACC; ACC = i + 1 

      7  => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC
      
      8  => "1111" & "000" & "001" & "000000000",  -- MOV ACC, R1
      
      9  => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC; ACC = ACC - R2
      10 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      -- 03: ST ACC,ACC  ; RAM[ACC] = ACC
      -- (endere�o = ACC, dado = ACC, coerente com sua liga��o RAM)
      11 => "0011" & "000" & "000" & "000000000",
      12 => "1010" & "011" & "000" & "000000000",  -- SUB, R3, ACC; ativar a flag negative
      13 => "0101" & "011" & "000" & "000000100",  -- BLT, R2, ACC, end4
      
      14 => "0000" & "000" & "000" & "000000000",
      
      ---- *****PASSO 2: eliminar os multiplos de 2, 3, 5 ****** ----
      ---- ***** eliminar multiplos de 2
      15 => "1001" & "000" & "000" & "000000010",  -- LD ACC, 2
      16 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      17 => "1001" & "000" & "000" & "000000010",
      18 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      19 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      20 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      21 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      22 => "1001" & "000" & "000" & "000100000",  -- LD ADD, 32
      23 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      24 => "0101" & "010" & "000" & "000010001",  -- BLT R2, ACC; end 17

      ---- ***** eliminar multiplos de 3
      25 => "1001" & "000" & "000" & "000000011",  -- LD ACC, 3
      26 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      27 => "1001" & "000" & "000" & "000000011",
      28 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      29 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      30 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      31 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      32 => "1001" & "000" & "000" & "000100000",  -- LD ADD, 32
      33 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      34 => "0101" & "010" & "000" & "000011011",  -- BLT R2, ACC; end 27

      ---- ***** eliminar multiplos de 5
      35 => "1001" & "000" & "000" & "000000101",  -- LD ACC, 5
      36 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      37 => "1001" & "000" & "000" & "000000101",
      38 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      39 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      40 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      41 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      42 => "1001" & "000" & "000" & "000100000",  -- LD ADD, 32
      43 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      44 => "0101" & "010" & "000" & "000100101",  -- BLT R2, ACC; end 37

      ---- ***** eliminar multiplos de 7
      45 => "1001" & "000" & "000" & "000000111",  -- LD ACC, 7
      46 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      47 => "1001" & "000" & "000" & "000000111",
      48 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      49 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      50 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      51 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      52 => "1001" & "000" & "000" & "000100000",  -- LD ADD, 32
      53 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      54 => "0101" & "010" & "000" & "000101111",  -- BLT R2, ACC; 47

      ---- ***** eliminar multiplos de 11
      55 => "1001" & "000" & "000" & "000001011",  -- LD ACC, 11
      56 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      57 => "1001" & "000" & "000" & "000001011",
      58 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      59 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      60 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      61 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      62 => "1001" & "000" & "000" & "000100000",  -- LD ADD, 32
      63 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      64 => "0101" & "010" & "000" & "000111001",  -- BLT R2, ACC; 57

      ---- *****PASSO 3: LOOP FINAL ****** ----
      65 => "1001" & "000" & "000" & "100000001",  -- LD ACC,#1
      
      66 => "1111" & "001" & "000" & "000000001",  -- MOV R1,ACC

      67 => "1001" & "000" & "000" & "000100000",  -- ACC = 32
      
      68 => "1111" & "010" & "000" & "000000000",  -- R2 = 32
      
      -- INICIO DO LOOP
      69 => "1001" & "000" & "000" & "000000000",  -- ACC = 0

      70 => "1111" & "011" & "000" & "000000000",  -- MOV, R3, ACC

      71 => "0110" & "001" & "000" & "000000000",  -- ADD, R1, ACC; ACC = i + 1 

      72 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC

      73 => "1111" & "000" & "001" & "000000000",  -- MOV ACC, R1
      
      74 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC; ACC = ACC - R2
      75 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      76 => "1010" & "011" & "000" & "000000000",  -- SUB, R3, ACC; ativar a flag negative
      77 => "0101" & "011" & "000" & "001000101",  -- BLT, R2, ACC, end69
      78 => "1001" & "000" & "000" & "000000001",  -- LD, ACC, 1
      79 => "1111" & "101" & "000" & "000000000",  -- MOV, R6, ACC
      80 => "0001" & "000" & "000" & "000000000",

      others => (others => '0')
   );
begin
   dado <= conteudo_rom(to_integer(endereco));
end architecture;