library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      endereco : in  unsigned(7 downto 0);
      dado     : out unsigned(18 downto 0)
   );
end entity;

architecture a_rom of rom is
   type mem is array (0 to 255) of unsigned(18 downto 0);

   constant conteudo_rom : mem := (
      ---- *****PASSO 1: colocar os valores de 1 a 32 ****** ----

      ---- SETUP INICIAL ----
      0  => "1001" & "000" & "000" & "000000001",  -- LD ACC,#1
      
      1  => "1111" & "001" & "000" & "000000001",  -- MOV R1,ACC

      2  => "1001" & "000" & "001" & "001100101",  -- ACC = 613
      
      3  => "1111" & "010" & "000" & "000000000",  -- R2 = 613
      
      -- INICIO DO LOOP
      4  => "1001" & "000" & "000" & "000000000",  -- ACC = 0

      5  => "1111" & "011" & "000" & "000000000",  -- MOV, R3, ACC

      6  => "0110" & "001" & "000" & "000000000",  -- ADD, R1, ACC; ACC = i + 1 

      7  => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC
      
      8  => "1111" & "000" & "001" & "000000000",  -- MOV ACC, R1
      
      9  => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC; ACC = ACC - R2
      10 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      -- 03: ST ACC,ACC  ; RAM[ACC] = ACC
      11 => "0011" & "000" & "000" & "000000000",
      12 => "1010" & "011" & "000" & "000000000",  -- SUB, R3, ACC; ativar a flag negative
      13 => "0101" & "011" & "000" & "000000100",  -- BLT, R3, ACC, end4
      
      14 => "0000" & "000" & "000" & "000000000",
      
      ---- *****PASSO 2: eliminar os multiplos de 2, 3, 5 ****** ----
      ---- ***** eliminar multiplos de 2
      15 => "1001" & "000" & "000" & "000000010",  -- LD ACC, 2
      16 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      17 => "1001" & "000" & "000" & "000000010",
      18 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      19 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      20 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      21 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      22 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      23 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      24 => "0101" & "010" & "000" & "000010001",  -- BLT R2, ACC; end 17

      ---- ***** eliminar multiplos de 3
      25 => "1001" & "000" & "000" & "000000011",  -- LD ACC, 3
      26 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      27 => "1001" & "000" & "000" & "000000011",
      28 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      29 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      30 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      31 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      32 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      33 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      34 => "0101" & "010" & "000" & "000011011",  -- BLT R2, ACC; end 27

      ---- ***** eliminar multiplos de 5
      35 => "1001" & "000" & "000" & "000000101",  -- LD ACC, 5
      36 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      37 => "1001" & "000" & "000" & "000000101",
      38 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      39 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      40 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      41 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      42 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      43 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      44 => "0101" & "010" & "000" & "000100101",  -- BLT R2, ACC; end 37

      ---- ***** eliminar multiplos de 7
      45 => "1001" & "000" & "000" & "000000111",  -- LD ACC, 7
      46 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      47 => "1001" & "000" & "000" & "000000111",
      48 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      49 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      50 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      51 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      52 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      53 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      54 => "0101" & "010" & "000" & "000101111",  -- BLT R2, ACC; 47

      ---- ***** eliminar multiplos de 11
      55 => "1001" & "000" & "000" & "000001011",  -- LD ACC, 11
      56 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      57 => "1001" & "000" & "000" & "000001011",
      58 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      59 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      60 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      61 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      62 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      63 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      64 => "0101" & "010" & "000" & "000111001",  -- BLT R2, ACC; 57
---- ***** eliminar multiplos de 13
      65 => "1001" & "000" & "000" & "000001101",  -- LD ACC, 13
      66 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      67 => "1001" & "000" & "000" & "000001101",  -- LD ACC, 13
      68 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      69 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      70 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      71 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      72 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      73 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      74 => "0101" & "010" & "000" & "001000011",  -- BLT R2, ACC; 67

      ---- ***** eliminar multiplos de 17
      75 => "1001" & "000" & "000" & "000010001",  -- LD ACC, 17
      76 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      77 => "1001" & "000" & "000" & "000010001",  -- LD ACC, 17
      78 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      79 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      80 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      81 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      82 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      83 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      84 => "0101" & "010" & "000" & "001001101",  -- BLT R2, ACC; 77

      ---- ***** eliminar multiplos de 19
      85 => "1001" & "000" & "000" & "000010011",  -- LD ACC, 19
      86 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      87 => "1001" & "000" & "000" & "000010011",  -- LD ACC, 19
      88 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      89 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      90 => "0011" & "000" & "011" & "000000000",  -- ST ACC, R3; RAM[ACC] = R3 = 0
      91 => "1111" & "010" & "000" & "000000000",  -- MOV, R2, ACC
      92 => "1001" & "000" & "001" & "001100101",  -- LD ADD, 613
      93 => "1010" & "010" & "000" & "000000000",  -- SUB R2, ACC
      94 => "0101" & "010" & "000" & "001011011",  -- BLT R2, ACC; 87

      ---- ***** eliminar multiplos de 23
      95 => "1001" & "000" & "000" & "000010111",  -- LD ACC, 23
      96 => "1111" & "001" & "000" & "000000000",  -- MOV R1, ACC
      -- INICIO DO LOOP
      97 => "1001" & "000" & "000" & "000010111",  -- LD ACC, 23
      98 => "0110" & "001" & "000" & "000000000",  -- ADD R1, ACC;
      99 => "1111" & "001" & "000" & "000000000",  -- MOV, R1, ACC;
      100 => "0011" & "000" & "011" & "000000000", -- ST ACC, R3; RAM[ACC] = R3 = 0
      101 => "1111" & "010" & "000" & "000000000", -- MOV, R2, ACC
      102 => "1001" & "000" & "001" & "001100101", -- LD ADD, 613
      103 => "1010" & "010" & "000" & "000000000", -- SUB R2, ACC
      104 => "0101" & "010" & "000" & "001100001", -- BLT R2, ACC; 97

      ---- *****PASSO 3: LOOP FINAL ****** ----
      105 => "1001" & "000" & "000" & "000000001", -- LD ACC,#1
      
      106 => "1111" & "001" & "000" & "000000001", -- MOV R1,ACC

      107 => "1001" & "000" & "001" & "001100101", -- ACC = 613
      
      108 => "1111" & "010" & "000" & "000000000", -- R2 = 613
      
      -- INICIO DO LOOP
      109 => "1001" & "000" & "000" & "000000000", -- ACC = 0

      110 => "1111" & "011" & "000" & "000000000", -- MOV, R3, ACC

      111 => "0110" & "001" & "000" & "000000000", -- ADD, R1, ACC; ACC = i + 1 

      112 => "1111" & "001" & "000" & "000000000", -- MOV, R1, ACC

      113 => "1111" & "000" & "001" & "000000000", -- MOV ACC, R1
      
      114 => "1010" & "010" & "000" & "000000000", -- SUB R2, ACC; ACC = ACC - R2
      115 => "1111" & "010" & "000" & "000000000", -- MOV, R2, ACC
      116 => "1010" & "011" & "000" & "000000000", -- SUB, R3, ACC; ativar a flag negative
      117 => "0101" & "011" & "000" & "001101101", -- BLT, R2, ACC, end109

      118 => "1001" & "000" & "000" & "101011111", -- LD ACC, RAM[607]
      119 => "0101" & "100" & "000" & "001111001", -- BLT R4, ACC (R4 = 0 por padrao), end122
      
      120 => "1001" & "000" & "000" & "000000001", -- LD ACC, 1
      121 => "1111" & "101" & "000" & "000000000", -- MOV, R5, ACC (R5 como bit debug)

      122 => "1001" & "000" & "000" & "000011111", -- LD, ACC, 31 (forcando ctz5)
      123 => "0110" & "101" & "000" & "000000000", -- ADD, R5, ACC (31 + 1)
      124 => "0010" & "000" & "000" & "001111110", -- CTZ5 126
      125 => "0000" & "000" & "000" & "000000000", -- NOP
      126 => "0001" & "000" & "000" & "000000000", -- HALT

      others => (others => '0')
   );
begin
   dado <= conteudo_rom(to_integer(endereco));
end architecture;