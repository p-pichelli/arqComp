library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      endereco : in  unsigned(7 downto 0);
      dado     : out unsigned(18 downto 0)
   );
end entity;

architecture a_rom of rom is
   type mem is array (0 to 255) of unsigned(18 downto 0);
   constant conteudo_rom : mem := (
      0 => "1001" & "000" & "000" & "100000101",  -- LD, imm=1, valor=5
      1 => "1111" & "011" & "000" & "000000000",  -- MOV R3 ? ACC
      
      2 => "1001" & "000" & "000" & "100001000",  -- LD, imm=1, val=8
      3 => "1111" & "100" & "000" & "000000000",  -- MOV R4? ACC
      4 => "0110" & "101" & "100" & "000000000",  -- ADD R5, src=R4
      5 => "1010" & "101" & "001" & "000000000",  -- SUB R5, src=R1
      6 => "1110" & "000" & "000" & "000010100", -- JUMP addr=20

      -- 7 => "1001" & "000" & "000" & "100000001",  -- LD, val=1
      -- 8 => "1111" & "001" & "000" & "000000000",  -- MOV R1 ? ACC
      -- 9 => "1111" & "000" & "101" & "000000000",  -- MOV ACC ? R5
      -- 10 => "1010" & "101" & "001" & "000000000",  -- SUB R5, src=R1
      7 => "1001" & "000" & "000" & "100000000",
      8 => "1111" & "101" & "000" & "000000000",
      9 => "0000000000000000000",
      10 => "0000000000000000000",
      11 => "0000000000000000000",
      12 => "0000000000000000000",
      13 => "0000000000000000000",
      14 => "0000000000000000000",
      15 => "0000000000000000000",
      16 => "0000000000000000000",
      17 => "0000000000000000000",
      18 => "0000000000000000000",
      19 => "0000000000000000000",
      20 => "1111" & "000" & "101" & "000000000", -- MOV ACC ?R5
      21 => "1111" & "011" & "000" & "000000000", -- MOV R3? ACC
      
      22 => "1110" & "000" & "000" & "000000100", -- JUMP addr=4
      
      23 => "1001" & "000" & "000" & "100000000",
      24 => "1111" & "011" & "000" & "000000000",
      
      others => "0000000000000000000"
   );
begin
   dado <= conteudo_rom(to_integer(endereco));
end architecture;
