library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      endereco : in  unsigned(7 downto 0);
      dado     : out unsigned(18 downto 0)
   );
end entity;

architecture a_rom of rom is
   type mem is array (0 to 255) of unsigned(18 downto 0);
   constant conteudo_rom : mem := (
      0 => "1001111000000000101",
      1 => "1111011111000000000",
      2 => "1001111000000001000",
      3 => "1111100111000000000",
      4 => "1111111011000000000",
      5 => "0110111100000000000",
      6 => "1111101111000000000",
      7 => "1001111000000000001",
      8 => "1010101111000000000",
      9 => "1110000000000010100",
      10 => "1001111000000000000",
      11 => "1111101111000000000",
      12 => "0000000000000000000",
      13 => "0000000000000000000",
      14 => "0000000000000000000",
      15 => "0000000000000000000",
      16 => "0000000000000000000",
      17 => "0000000000000000000",
      18 => "0000000000000000000",
      19 => "0000000000000000000",
      20 => "1111111101000000000",
      21 => "1111011111000000000",
      22 => "1110000000000000100",
      23 => "1001111000000000000",
      24 => "1111011111000000000",
      others => "0000000000000000000"
   );
begin
   dado <= conteudo_rom(to_integer(endereco));
end architecture;
