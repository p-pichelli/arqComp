library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      endereco : in  unsigned(7 downto 0);
      dado     : out unsigned(18 downto 0)
   );
end entity;

architecture a_rom of rom is
   type mem is array (0 to 255) of unsigned(18 downto 0);
   constant conteudo_rom : mem := (
      0  => "000000000000000000000001", -- LW mem�ria[1]
      1  => "000000000000000000000010", -- LW mem�ria[2]
      2  => "000100000000000000000000", -- ADD R0
      3  => "000100000001000000000000", -- ADD R1
      4  => "001000000010000000000000", -- SUB R2
      5  => "001000000011000000000000", -- SUB R3
      6  => "010000000100000000000000", -- AND R4
      7  => "010000000101000000000000", -- AND R5
      8  => "010100000000000000000000", -- OR R0
      9  => "010100000001000000000000", -- OR R1
      10 => "001100000000000000000011", -- SW mem�ria[3]
      11 => "001100000000000000000100", -- SW mem�ria[4]
      12 => "011100000000000000001100", -- BR se acumulador=0 ROM[12]
      13 => "100000000000000000010100", -- JMP ROM[20]
      14 => "111100000000000000000000", -- NOP
      15 => "000000000000000000000101", -- LW mem�ria[5]
      16 => "000100000010000000000000", -- ADD R2
      17 => "001000000011000000000000", -- SUB R3
      18 => "010000000001000000000000", -- AND R1
      19 => "010100000100000000000000", -- OR R4
      20 => "001100000000000000000101", -- SW mem�ria[5]
      21 => "011100000000000000010101", -- BR se acumulador=0 ROM[21]
      22 => "100000000000000000011000", -- JMP ROM[24]
      23 => "111100000000000000000000", -- NOP
      24 => "000000000000000000000110", -- LW mem�ria[6]
      25 => "000100000011000000000000", -- ADD R3
      26 => "001000000100000000000000", -- SUB R4
      27 => "010000000101000000000000", -- AND R5
      28 => "010100000010000000000000", -- OR R2
      29 => "001100000000000000000110", -- SW mem�ria[6]
      30 => "011100000000000000011110", -- BR se acumulador=0 ROM[30]
      31 => "100000000000000000100000", -- JMP ROM[32]
      32 => "111100000000000000000000", -- NOP
      33 => "000000000000000000000111", -- LW mem�ria[7]
      34 => "000100000001000000000000", -- ADD R1
      35 => "001000000010000000000000", -- SUB R2
      36 => "010000000011000000000000", -- AND R3
      37 => "010100000100000000000000", -- OR R4
      38 => "001100000000000000000111", -- SW mem�ria[7]
      39 => "011100000000000000101000", -- BR se acumulador=0 ROM[40]
      40 => "100000000000000000101000", -- JMP ROM[40]
      41 => "111100000000000000000000", -- NOP
      42 => "000000000000000000001000", -- LW mem�ria[8]
      43 => "000100000010000000000000", -- ADD R2
      44 => "001000000011000000000000", -- SUB R3
      45 => "010000000001000000000000", -- AND R1
      46 => "010100000100000000000000", -- OR R4
      47 => "001100000000000000001000", -- SW mem�ria[8]
      48 => "011100000000000000110010", -- BR se acumulador=0 ROM[50]
      49 => "100000000000000000110010", -- JMP ROM[50]
      others => "111100000000000000000000" -- NOP
   );
begin
   dado <= conteudo_rom(to_integer(endereco));
end architecture;
